/*========================================================
File name:      defines.sv
Description:    APB defines file
Author:         Jaimil Patel
Date created:   21 June 2020
=========================================================*/

`define TOTAL_NUMBER_OF_SLAVES 8'd1

`define APB_REG_ADDR_HIGH 31
`define APB_REG_ADDR_LOW  0

`define APB_REG_DATA_HIGH 31
`define APB_REG_DATA_LOW  0

`define APB_REG_STROBE_HIGH 7
`define APB_REG_STROBE_LOW  0


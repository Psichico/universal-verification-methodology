/*========================================================
File name:      interface.sv
Description:    template
Author:         Jaimil Patel
Date created:   18 June 2020
=========================================================*/

interface interface_template(input logic clock);

    //logic [7:0] a;
    //logic [7:0] b;

endinterface: interface_template

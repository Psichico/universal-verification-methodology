/*========================================================
File name:      interface.sv
Description:    APB interface
Author:         Jaimil Patel
Date created:   21 June 2020
=========================================================*/

interface apb_interface(input logic clock);


endinterface: apb_interface
